library verilog;
use verilog.vl_types.all;
entity group32_hw5_vlg_vec_tst is
end group32_hw5_vlg_vec_tst;
