library verilog;
use verilog.vl_types.all;
entity group32_hw6_vlg_vec_tst is
end group32_hw6_vlg_vec_tst;
